library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity clkDiv is
   port(  clk100, Reset: in std_logic; -- Entrees du diviseur d'horloge
          clk25:         out std_logic); --Horloge de sortie
end clkDiv;

architecture divHorl of clkDiv is
    
signal compt: std_logic_vector(1 downto 0); -- compteur

begin
    
	-- Gestion du diviseur d'horloge
    process (clk100,Reset)
    begin
    	if (Reset='0') then compt<="00";
	elsif rising_edge(clk100) then compt<=compt+'1';
	end if;
    end process;
    
    clk25<=compt(1);

end divHorl;